module instruction_memory(output[31:0] instruction, input[31:0] read_instruct_addr);
reg[7:0] mem[0:255];
initial begin
	 $readmemb("instruction_list.txt", mem);
			 
			 /* mem[0]=32'b100011_11101_00001_0000000000000000
				mem[4]=32'b100011_11101_00010_0000000000000001
				mem[8]=32'b100011_11101_00011_0000000000000010
				mem[12]=32'b100011_11101_00000_0000000000000000
				mem[16]=32'b100011_11101_00101_0000000000000000
				mem[20]=32'b100011_11101_00110_0000000000000011
				mem[24]=32'b100011_11101_00111_0000000000000100

				mem[28]=32'b000101_00001_00000_0000000000001101.....13 or 14....32
				mem[32]=32'b000000_00010_00011_00100_00000_101011
				mem[36]=32'b000101_00100_00000_0000000000000011	...3 or 4...line40
				mem[40]=32'b000101_00011_00000_0000000000001000....10 or 11...line44
				mem[44]=32'b000000_00001_00110_00001_00000_100101
				mem[48]=32'b000010_1111_1111_1111_1111_1111_11_1010			.........j -6
				000000_00101_00000_00101_100100
				mem[52]=32'b000000_00101_00010_00101_00000_100101
				mem[56]=32'b000000_00010_00000_00010_00000_100100
				mem[60]=32'b000000_00010_00011_00010_00000_100101
				mem[64]=32'b000000_00011_00000_00011_00000_100100
				mem[68]=32'b000000_00011_00101_00011_00000_100101
				mem[72]=32'b000010_1111_1111_1111_1111_1111_11_0100			........j -12

				mem[76]=32'b000000_00010_00011_00010_00000_100010
				mem[80]=32'b000010_1111_1111_1111_1111_1111_11_0010			......j -14

				mem[84]=32'b000000_00111_00010_00111_00000_100101
				mem[88]=32'b101011_11101_00111_0000000000000100
				mem[89]=32'b000010_1111_1111_1111_1111_1111_11_0001	
		*/



end


assign	instruction ={mem[read_instruct_addr],
				   mem[read_instruct_addr+1],
				   mem[read_instruct_addr+2],
				   mem[read_instruct_addr+3]};

endmodule
